`define subFrameH 64
`define subFrameV 64
`define overlapH 32
`define overlapV 32
`define rangeH 7
`define rangeV 7
`define possibleH `rangeH * `overlapH //32*7
`define possibleV `rangeV * `overlapV //32*7

`define gradeFactor 5
