//**************************************
// File Name        : Top.sv
// Created Time     : 2025/05/15 20:00
// Last Revised Time: 2025/05/15 21:00
//**************************************

module Top (
  input i_clk,
  input i_rst_n
);
  
endmodule